module adder (
    input  [14:0] a,
    b,
    output [14:0] y
);
  assign y = a + b;
endmodule
