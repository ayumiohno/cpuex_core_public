module adder (
    input  [17:0] a,
    b,
    output [17:0] y
);
  assign y = a + b;
endmodule
